`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name: SevenSegmentDisplay
// Description: 
//////////////////////////////////////////////////////////////////////////////////


module SevenSegmentDisplay(

    );
endmodule
